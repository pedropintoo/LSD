-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.1 Build 720 11/11/2020 SJ Lite Edition
-- Created on Thu Apr 06 12:49:46 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

ENTITY DrinksFSM IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        V : IN STD_LOGIC := '0';
        C : IN STD_LOGIC := '0';
        abrir : OUT STD_LOGIC;
		  currentState : out std_logic_vector(3 downto 0)
    );
END DrinksFSM;

ARCHITECTURE BEHAVIOR OF DrinksFSM IS
    TYPE type_fstate IS (E0,E1,E2,E3,E4,E5);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,V,C)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= E0;
            abrir <= '0';
        ELSE
            abrir <= '0';
            CASE fstate IS
                WHEN E0 =>
                    IF ((NOT((C = '1')) AND (V = '1'))) THEN
                        reg_fstate <= E1;
                    ELSIF ((C = '1')) THEN
                        reg_fstate <= E3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E0;
                    END IF;

                    abrir <= '0';
                WHEN E1 =>
                    IF ((NOT((C = '1')) AND (V = '1'))) THEN
                        reg_fstate <= E2;
                    ELSIF ((C = '1')) THEN
                        reg_fstate <= E4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E1;
                    END IF;

                    abrir <= '0';
                WHEN E2 =>
                    IF ((NOT((C = '1')) AND (V = '1'))) THEN
                        reg_fstate <= E3;
                    ELSIF ((C = '1')) THEN
                        reg_fstate <= E5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E2;
                    END IF;

                    abrir <= '0';
                WHEN E3 =>
                    IF ((NOT((C = '1')) AND (V = '1'))) THEN
                        reg_fstate <= E4;
                    ELSIF ((C = '1')) THEN
                        reg_fstate <= E5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E3;
                    END IF;

                    abrir <= '0';
                WHEN E4 =>
                    IF (((V = '1') OR (C = '1'))) THEN
                        reg_fstate <= E5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E4;
                    END IF;

                    abrir <= '0';
                WHEN E5 =>
                    reg_fstate <= E0;

                    abrir <= '1';
                WHEN OTHERS => 
                    abrir <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
	 
	 					
	-- converts an enumerated type type_fstate into a 4-bit std_logic_vector.	
	currentState <= std_logic_vector(to_unsigned(type_fstate'pos(reg_fstate),4));
	
END BEHAVIOR;
